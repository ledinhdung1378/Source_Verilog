module tb_register_4bit ;

reg clk,clr,ce ; 
reg d[3:0] ; 
wire q[3:0] ; 

register_4bit uut (.clk(clk),.clr(clr),.d(d),.q(q)) ; 

initial    
    begin 
        clr = 0 ; 
        forever #5 clk = ~clk ; 
    end 

initial 
    begin 
        clr = 0 ;
        ce = 0 ;
        d = 4'b1011 ; 
        #10 ; 
        ce = 1 ; 
        d = 4'b1000 ; 
        #10 ;
        d = 4'b0001 ; 
        #10 ; 
        clr = 1; 
        #10 ; 
        clr = 0 ; 
        d = 4'b1111; 
        #10 ; 
        $finish ; 
    end 

endmodule ;     